
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE WORK.PACK.ALL;

entity COM_BUS is
	PORT(
		S: IN STD_LOGIC_VECTOR(3 DOWNTO 0); --SELECT LINES
		-- BUS OUTPUT
		DATA_BUS_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		-- BUS INPUTS
		DATA_AR : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		DATA_PC : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		DATA_DR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		DATA_AC : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		DATA_IR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		DATA_MEM : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
                DATA_TR : IN STD_LOGIC_VECTOR(15 DOWNTO 0); 
          
	);
end COM_BUS;

architecture Behavioral of COM_BUS is
SIGNAL DATA_NULL : STD_LOGIC_VECTOR (7 DOWNTO 0):=(OTHERS=>'Z');
begin
	-- TAKES ALL INPUTS
	-- RETURNS OUTPUT IN DATA_BUS_OUT
	MUX : MUX8X1_V8 PORT MAP (DATA_PC,DATA_AR,DATA_DR,DATA_AC,DATA_MEM,DATA_IR, DATA_TR, DATA_NULL, S, DATA_BUS_OUT);    
	
end Behavioral;
